module maindec(input    logic [6:0] op,
                           output logic [1:0] ResultSrc,
                           output logic           MemWrite,
                           output logic           Branch, ALUSrc,
                           output logic           RegWrite, Jump,
                           output logic [1:0] ImmSrc,
                           output logic [1:0] ALUOp,
                           output logic           RegWrite_for_hazard
                           );
    logic [10:0] controls;
    logic RegWrite_for_hazard;
    assign {RegWrite_s, ImmSrc_s, ALUSrc_s, MemWrite_s,
                  ResultSrc_s, Branch_s, ALUOp_s, Jump_s} = controls;

      signal_history #(  
      .WIDTH(2),
      .DEPTH(3)
      ) result_src_reg(
      clk,
      reset,
      ResultSrc_s,
      ResultSrc
   );
   flopr #(32) last_flop_for_regwrite (
      clk,
      reset,
      RegWrite_for_hazard,
      RegWrite
   );

   signal_history #(    
      .WIDTH(1),
      .DEPTH(2)
    ) register_write_reg(
      clk,
      reset,
      RegWrite_s,
      RegWrite_for_hazard
   );
   signal_history #(  
      .WIDTH(1),
      .DEPTH(2)
      ) mem_write_reg(
      clk,
      reset,
      MemWrite_s,
      MemWrite
   );
   //delay ALU_src only 1 clock
   flopr #(32) pcreg (
      clk,
      reset,
      ALUSrc_s,
      ALUSrc
   );
   //delay jump_S only 1 clock
   flopr #(32) pcreg (
      clk,
      reset,
      Jump_s,
      Jump
   );
   //delay branchD only 1 clock
   flopr #(32) pcreg (
      clk,
      reset,
      Branch_s,
      Branch
   );

    always_comb
       case(op)
       // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
            7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
          7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
          7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type
          7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
          7'b0010011: controls = 11'b1_00_1_0_00_0_10_0; // I-type ALU
          7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal
           default:      controls = 11'bx_xx_x_x_xx_x_xx_x; // ??? 
        endcase
endmodule