//*Suman 2 del reg 1 al 12

00200093//ADDI x1, x0, 1
00200113//ADDI x2, x0, 2
00200193//ADDI x3, x0, 3
00200213//ADDI x4, x0, 4
00200313//ADDI x5, x0, 5
00200393//ADDI x6, x0, 6
00200413//ADDI x7, x0, 7
00200493//ADDI x8, x0, 8
00200513//ADDI x9, x0, 9
00200593//ADDI x10, x0, 10
00200613//ADDI x11, x0, 11

///////////111///////

01400093 //* addi x10, x1, 20 


/////////////////

00000093 //ADDI x1, x0, 0
00000113 //ADDI x2, x0, 0
00000193 //ADDI x3, x0, 0
00000213 //ADDI x4, x0, 0
00000293 //ADDI x5, x0, 0
00000313 //ADDI x6, x0, 0
00000393 //ADDI x7, x0, 0
00000413 //ADDI x8, x0, 0
00000493 //ADDI x9, x0, 0
00000513 //ADDI x10, x0, 0
00000593 //ADDI x11, x0, 0
00000613 //ADDI x12, x0, 0
00000693 //ADDI x13, x0, 0
00000713 //ADDI x14, x0, 0
00000793 //ADDI x15, x0, 0
00000813 //ADDI x16, x0, 0
00000893 //ADDI x17, x0, 0
00000913 //ADDI x18, x0, 0
00000993 //ADDI x19, x0, 0
00000A13 //ADDI x20, x0, 0
00000A93 //ADDI x21, x0, 0
00000B13 //ADDI x22, x0, 0
00000B93 //ADDI x23, x0, 0
00000C13 //ADDI x24, x0, 0
00000C93 //ADDI x25, x0, 0
00000D13 //ADDI x26, x0, 0
00000D93 //ADDI x27, x0, 0
00000E13 //ADDI x28, x0, 0
00000E93 //ADDI x29, x0, 0
00000F13 //ADDI x30, x0, 0
00000F93 //ADDI x31, x0, 0

//*AND I
00210593   // andi x11, x2, 2
00310613   // andi x12, x3, 3
00410693   // andi x13, x4, 4
00510713   // andi x14, x5, 5
00610793   // andi x15, x6, 6
//*ORI
00710813   // ori x16, x7, 7
00810893   // ori x17, x8, 8
00910913   // ori x18, x9, 9
00A10993   // ori x19, x10, 10
//*
0023E2B3  // or x7,  x7, x2    # x7 = (x7 OR x2)
0023E3B3 // or x8,  x7, x2    # x8 = (x7 OR x2)
0023E4B3 // or x9,  x7, x2    # x9 = (x7 OR x2)
0023E5B3 // or x10, x7, x2    # x10 = (x7 OR x2)
00326BB3 // or x23, x4, x3    # x23 = (x4 OR x3)
00326C33 // or x24, x4, x3    # x24 = (x4 OR x3)
00326CB3 // or x25, x4, x3    # x25 = (x4 OR x3)
00326D33 // or x26, x4, x3    # x26 = (x4 OR x3)
00326DB3 // or x27, x4, x3    # x27 = (x4 OR x3)
00326E33 // or x28, x4, x3    # x28 = (x4 OR x3)
00326EB3 // or x29, x4, x3    # x29 = (x4 OR x3)
00326F33 // or x30, x4, x3    # x30 = (x4 OR x3)





















//!---------------------------No andan por bug del rd = al inmediatio que no tiene sentido
00100093 // addi x1, x0, 1
00200113 // addi x2, x0, 2
00300193 // addi x3, x0, 3
00400213 // addi x4, x0, 4
00500293 // addi x5, x0, 5
00600313 // addi x6, x0, 6
00700393 // addi x7, x0, 7
00800413 // addi x8, x0, 8
00900493 // addi x9, x0, 9
00A00513 // addi x10, x0, 10
00B00593 // addi x11, x0, 11
00C00613 // addi x12, x0, 12
00D00693 // addi x13, x0, 13
00E00713 // addi x14, x0, 14
00F00793 // addi x15, x0, 15
01000813 // addi x16, x0, 16
01100893 // addi x17, x0, 17
01200913 // addi x18, x0, 18
01300993 // addi x19, x0, 19
01400A13 // addi x20, x0, 20
01500A93 // addi x21, x0, 21
01600B13 // addi x22, x0, 22
01700B93 // addi x23, x0, 23
01800C13 // addi x24, x0, 24
01900C93 // addi x25, x0, 25
01A00D13 // addi x26, x0, 26
01B00D93 // addi x27, x0, 27
01C00E13 // addi x28, x0, 28
01D00E93 // addi x29, x0, 29
01E00F13 // addi x30, x0, 30
01F00F93 // addi x31, x0, 31
///////////////////////